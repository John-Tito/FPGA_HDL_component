//---------------------------------------------------------------------------------------
// uart transmit module
//
//---------------------------------------------------------------------------------------
// verilog_format: off
`resetall
`timescale 1ns / 1ps
`default_nettype none
// verilog_format: on
module uart_tx (
    input  wire       clock,        // global clock input
    input  wire       reset,        // global reset input
    input  wire       ce_16,        // baud rate multiplyed by 16 - generated by baud module
    input  wire [7:0] tx_data,      // data byte to transmit
    input  wire       tx_new_data,  // asserted to indicate that there is a new data byte for transmission
    input  wire       send_parity,  // asserted to indicate that there is a parity bit
    input  wire       odd_even,     // asserted to indicate that the parity bit is odd or even
    output reg        ser_out,      // serial data output
    output reg        tx_busy       // signs that transmitter is busy
);
    //---------------------------------------------------------------------------------------
    // modules inputs and outputs


    // internal wires
    wire ce_1;  // clock enable at bit rate

    wire [3:0] data_length;

    // internal registers
    reg [3:0] count16;
    reg [3:0] bit_count;
    reg [8:0] data_buf;
    reg parity_bit;
    //---------------------------------------------------------------------------------------
    // module implementation
    // a counter to count 16 pulses of ce_16 to generate the ce_1 pulse
    always @(posedge clock or posedge reset) begin

        if (reset) count16 <= 4'b0;
        else if (tx_busy & ce_16) count16 <= count16 + 4'b1;
        else if (~tx_busy) count16 <= 4'b0;

    end

    // ce_1 pulse indicating output data bit should be updated
    assign ce_1        = (count16 == 4'b1111) & ce_16;

    assign data_length = (send_parity) ? 4'd10 : 4'd9;

    // tx_busy flag
    always @(posedge clock or posedge reset) begin
        if (reset) tx_busy <= 1'b0;
        else if (~tx_busy & tx_new_data) tx_busy <= 1'b1;
        else if (tx_busy & (bit_count == data_length) & ce_1) tx_busy <= 1'b0;
    end

    // output bit counter
    always @(posedge clock or posedge reset) begin
        if (reset) bit_count <= 4'h0;
        else if (tx_busy & ce_1) bit_count <= bit_count + 4'h1;
        else if (~tx_busy) bit_count <= 4'h0;
    end

    // data shift register
    always @(posedge clock or posedge reset) begin
        if (reset) begin
            data_buf   <= 9'b0;
            parity_bit <= 0;
        end else if (~tx_busy) begin
            data_buf   <= {tx_data, 1'b0};
            parity_bit <= 0;
        end else if (tx_busy & ce_1) begin
            if (send_parity) begin
                if (bit_count <= 4'd7) begin
                    data_buf   <= {1'b1, data_buf[8:1]};
                    parity_bit <= parity_bit + data_buf[1];
                end else if (bit_count == 4'd8) begin
                    if (odd_even) data_buf <= {data_buf[8:1], ~parity_bit};
                    else data_buf <= {data_buf[8:1], parity_bit};
                end else begin
                    data_buf <= {1'b1, data_buf[8:1]};
                end
            end else begin
                data_buf <= {1'b1, data_buf[8:1]};
            end
        end
    end

    // output data bit
    always @(posedge clock or posedge reset) begin
        if (reset) ser_out <= 1'b1;
        else if (tx_busy) ser_out <= data_buf[0];
        else ser_out <= 1'b1;
    end

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------
